//
// lab8 : version 06/12/2020
// 
`timescale 1ns/1ps


module sw_decode (output logic bits_done, output logic bit_value,
	input logic next_bit, input logic [10:0] sw,
	input logic clk, input logic rst);

	// enter your code here


endmodule
