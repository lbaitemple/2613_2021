//
// lab3 : version 06/12/2020
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module svn_seg_decoder(
	output logic [6:0] seg_out,
	input logic [3:0] bcd_in,
	input logic display_on
	);

	// add the design code here

endmodule
