module and_3_inputs (output logic f, input logic a, b, c);
	// this is the design to test
	assign f = a & b & c;
endmodule
