`timescale 1ns / 1ps

module up_down_count_dp (output logic [3:0] digit3, output logic [3:0] digit2,
	output logic [3:0] digit1, output logic [3:0] digit0,
	input logic enable, input logic up_down, input logic rst, input clk);

	logic c_out0, c_out1, c_out2;	// internal carry out signals

        // instantiate the 4 binary coded decimal counters

endmodule
