{"filter":false,"title":"tb_gates.sv","tooltip":"/lab1/tb_gates.sv","ace":{"folds":[],"scrolltop":312,"scrollleft":0,"selection":{"start":{"row":19,"column":16},"end":{"row":19,"column":16},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":0},"hash":"e7533ef4450a55c9e14114e9379fe3b9701fdb96","undoManager":{"mark":-1,"position":-1,"stack":[]},"timestamp":1534119608000}