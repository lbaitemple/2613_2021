//
// lab7 : version 01/04/20205
//  
`timescale 1ns/1ps

module ir_emitter_dp (output logic emitter_out, output logic tc_modulator, input logic clk,
	input logic rst, input logic ena, input [1:0] mod_sel, input logic sw_modulator);

	// enter your code here

endmodule
