{"filter":false,"title":"tb_memory_display.sv","tooltip":"/lab11/tb_memory_display.sv","undoManager":{"mark":-1,"position":-1,"stack":[]},"ace":{"folds":[],"scrolltop":1114.5,"scrollleft":1.5,"selection":{"start":{"row":0,"column":0},"end":{"row":0,"column":0},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":{"row":68,"state":"start","mode":"ace/mode/verilog"}},"timestamp":1592406716365,"hash":"c5e3e7194713d56f03c110d3798c71c91a09002a"}