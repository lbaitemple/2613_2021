//
// lab10 : version 03/29/2020
//  
`timescale 1ns/1ps

module ir_emitter_fsm (output logic sw_modulator, output logic [1:0] mod_sel, output logic dp_rst,
	output logic next_bit, input logic clk, input logic rst, input logic strt,
	input logic tc_modulator, input logic bits_done, input logic bit_value);

	// enter your code here

endmodule
