{"filter":false,"title":"hamming7_4_decode.sv","tooltip":"/lab4/hamming7_4_decode.sv","undoManager":{"mark":-1,"position":-1,"stack":[]},"ace":{"folds":[],"scrolltop":0,"scrollleft":0,"selection":{"start":{"row":0,"column":0},"end":{"row":0,"column":0},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":0},"timestamp":1592311614907,"hash":"69da6caf47ab6dfc7e41602d79fec5ed82c565e7"}