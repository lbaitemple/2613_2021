//
// lab2 : version 06/12/2020
// 
`timescale 1ns / 1ps
module hamming7_4_encode(
	output logic [7:1] e,
	input logic [4:1] d
	);

	// enter your code here

endmodule
