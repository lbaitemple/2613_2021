//
// lab8 : version 01/01/2025
// 

module memory_display (output logic [6:0] cathode, output logic [3:0] anode,
	input logic rst, input logic clk, 
	output logic [3:0] rs_data, output logic [3:0] ru_data,
	input logic w_ena, input logic [3:0] w_data, input logic [9:0] sw);



endmodule
