//
// lab6 : version 06/12/2020
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module alu_1 (output logic [3:0] f, output logic c_out, input logic [2:0] sel,
	input logic [3:0] a, input logic [3:0] b, input logic c_in);

	// enter your code here

endmodule
