//
// lab7 : version 01/04/2025
//  
module divider #(parameter BIT_SIZE=4)
	(output logic tc, output logic [BIT_SIZE-1:0] count, input logic clk,
	input logic rst, input logic ena, input logic [BIT_SIZE-1:0] init_count);

	// enter your code here


endmodule