`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module lab3_decoder(
	output logic [3:0] an,
	output logic [6:0] cathode,
	input logic [6:0] sw
	);

	// instantiate two outputs from the class presentation, double check with your TA for the values 
	assign an = [];
	assign cathode =[];

endmodule
