{"changed":false,"filter":false,"title":"tb_lab4_decoder.sv","tooltip":"/lab4/tb_lab4_decoder.sv","value":"`timescale 1ns / 1ps\n////////////////////////////////////////////////////////////////////////////////\n////////////////////////////////////////////////////////////////////////////////\n\nmodule tb_lab4_decoder;\n\n\t// Inputs\n\tlogic [6:0] h_code;\n\n\t// Outputs\n\tlogic [6:0] segment;\n\tlogic [3:0] data_out;\n\tlogic [3:0] an;\n\n\t// Instantiate the Unit Under Test (UUT)\n\tlab4_decoder uut (.led(data_out), .an, .cathode(segment), .sw(h_code));\n\t\n\t// parameters of test vectors (outputs = columns - inputs)\n\tparameter COLUMNS = 18, INPUTS = 7, ROWS = 128;\n\n\t// this is how you declare a two dimensional test vector\n\tlogic [COLUMNS-1:0] test_vector [0:ROWS-1];\n\t// we need a single vector also to make things easy\n\tlogic [COLUMNS-1:0] single_vector;\n\tinteger i;\t// and define a variable for an index\n\tinteger mm_count;\t// define a variable to count mismatches\n\n\tinitial begin\n\t\t$dumpfile(\"tb_lab4_decoder.vcd\");\n\t\t$dumpvars();\n\n\t\tmm_count = 0;\t// zero mismatch count\n\n\t\t// first read all of the test vectors from a file into array: test_vector\n\t\t$readmemb(\"tb_lab4_decoder.txt\", test_vector);\n\t\t\n\t\t// need to loop over all of the rows using a for loop\n\t\tfor (i=0; i<ROWS; i=i+1) begin\n\t\t\t// put the vector to test this loop into single_vector\n\t\t\tsingle_vector = test_vector [i];\n\t\t\t\n\t\t\t// now apply the stimuli to from the vector to the input signals\n\t\t\th_code = single_vector[COLUMNS-1:COLUMNS-INPUTS];\n\t\t\t#10;\t// wait 10 ns for inputs to settle\n\t\t\t// compare to expected value\n\t\t\tif ({segment,data_out} !== single_vector[COLUMNS-INPUTS-1:0]) begin\n\t\t\t\t// display mismatch\n\t\t\t\t$display(\"Mismatch--loop index i: %d; input: %b, expected: %b_%b, received: %b_%b\",\n\t\t\t\t\ti, h_code, single_vector[COLUMNS-INPUTS-1:4],\n\t\t\t\t\tsingle_vector[3:0], segment, data_out);\n\n\t\t\t\tmm_count = mm_count + 1;\t// increment mismatch count\n\n\t\t\tend\n\t\t\t#10;\t// add 10 ns for symmetry\n\t\tend\t// end of for loop\n\n\t\t// tell designer we're done with the simulation\n\t\tif (mm_count == 0) begin\n\t\t\t$display(\"Simulation complete - no mismatches!!!\");\n\t\tend else begin\n\t\t\t$display(\"Simulation complete - %d mismatches!!!\", mm_count);\n\t\tend\n\t\t$finish;\n\t\t\n\tend\t// end of initial block\nendmodule\n","undoManager":{"mark":-1,"position":-1,"stack":[]},"ace":{"folds":[],"scrolltop":0,"scrollleft":0,"selection":{"start":{"row":0,"column":0},"end":{"row":0,"column":0},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":0},"timestamp":1534122029000}