{"filter":false,"title":"tb_hamming7_4_decode.sv","tooltip":"/lab4/tb_hamming7_4_decode.sv","ace":{"folds":[],"scrolltop":382.5,"scrollleft":0,"selection":{"start":{"row":0,"column":0},"end":{"row":0,"column":0},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":0},"hash":"02746b7e259ad076306d82a3e9a811baaec411b4","undoManager":{"mark":-1,"position":-1,"stack":[]},"timestamp":1534121953000}