{"filter":false,"title":"gates.sv","tooltip":"/lab1/gates.sv","undoManager":{"mark":-1,"position":-1,"stack":[]},"ace":{"folds":[],"scrolltop":0,"scrollleft":0,"selection":{"start":{"row":13,"column":0},"end":{"row":13,"column":0},"isBackwards":false},"options":{"guessTabSize":true,"useWrapMode":false,"wrapToView":true},"firstLineState":{"row":24,"mode":"ace/mode/verilog"}},"timestamp":1591975277891,"hash":"93bd126a1cef9ceebccb13de5839fa53bb04f10e"}